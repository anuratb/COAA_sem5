`timescale 1ns / 1ps

////////////////////////////////////////////////////////////////////////////////
// Anurat Bhattacharya : 19CS10071
// Sunanda Mandal : 19CS10060
//
// Create Date:   11:14:47 08/25/2021
// Design Name:   RCA64
// Module Name:   /home/ise/COAA_Assign1/rca64_tb.v
// Project Name:  COAA_Assign1
// Target Device:  
// Tool versions:  
// Description: 
//
// Verilog Test Fixture created by ISE for module: RCA64
//
// Dependencies:
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
////////////////////////////////////////////////////////////////////////////////

module rca64_tb;

	// Inputs
	reg [63:0] A1;
	reg [63:0] A2;
	reg in;

	// Outputs
	wire [63:0] S;
	wire C;

	// Instantiate the Unit Under Test (UUT)
	RCA64 uut (
		.A1(A1), 
		.A2(A2), 
		.in(in), 
		.S(S), 
		.C(C)
	);

	initial begin
		// Initialize Inputs
		A1 = 0;
		A2 = 0;
		in = 0;

		// Wait 100 ns for global reset to finish
		#100;
		
        
		// Add stimulus here
		#2
		begin
			A1 = 64'b111000011000001110011101111101100110100001000000101010101101010;
			A2 = 64'b100100110000110110000011000111100101011011111101101010111;
			in = 1;
			$monitor("A1 = %b, A2 = %b,in = %b : S = %b,C=%b",A1,A2,in,S,C);
		end
		#2
		begin
			A1 = 64'b110111000010010100110101111001100111111011011111101110011000001;
			A2 = 64'b101110111001000111011000000101001001010101100100100110111101010;
			in = 0;
			$monitor("A1 = %b, A2 = %b,in = %b : S = %b,C=%b",A1,A2,in,S,C);
		end
		#2
		begin
			A1 = 64'b101100111111101100011110001101101111000011000001100010100000110;
			A2 = 64'b110110110101111100110011000010001001111010001101010110110111100;
			in = 1;
			$monitor("A1 = %b, A2 = %b,in = %b : S = %b,C=%b",A1,A2,in,S,C);
		end
		#2
		begin
			A1 = 64'b1101100011001011111011111001100110111100001011111110001000001;
			A2 = 64'b111110100110010111011000110011000110011110000001110111011010100;
			in = 1;
			$monitor("A1 = %b, A2 = %b,in = %b : S = %b,C=%b",A1,A2,in,S,C);
		end
		#2
		begin
			A1 = 64'b10001110010011011111111001010101110110111010000000111111100100;
			A2 = 64'b11100111010110001100111101101001101011110110100100001001011101;
			in = 1;
			$monitor("A1 = %b, A2 = %b,in = %b : S = %b,C=%b",A1,A2,in,S,C);
		end
		#2
		begin
			A1 = 64'b111010001110111101100000001010001010000011111000011011000101001;
			A2 = 64'b101100011011101000100010110110100111001000010001101000101000111;
			in = 1;
			$monitor("A1 = %b, A2 = %b,in = %b : S = %b,C=%b",A1,A2,in,S,C);
		end
		#2
		begin
			A1 = 64'b110110100101001001001101011000101010000011101010011001010101011;
			A2 = 64'b10100111010111001000100000100001010101110111100101001110010000;
			in = 0;
			$monitor("A1 = %b, A2 = %b,in = %b : S = %b,C=%b",A1,A2,in,S,C);
		end
		#2
		begin
			A1 = 64'b1010101001110001100000101000101001010110001001111101101101110;
			A2 = 64'b110000000000000011111100011101101101001100110100011000110111100;
			in = 1;
			$monitor("A1 = %b, A2 = %b,in = %b : S = %b,C=%b",A1,A2,in,S,C);
		end
		#2
		begin
			A1 = 64'b110000111111010111101101100001101110101101100101010100100000110;
			A2 = 64'b11000101000001101001000111111100000101001001001010000001010111;
			in = 0;
			$monitor("A1 = %b, A2 = %b,in = %b : S = %b,C=%b",A1,A2,in,S,C);
		end
		#2
		begin
			A1 = 64'b11110010101010100111001001100000100111101011011010011011011010;
			A2 = 64'b111000001101011100010110110110101111010110001010111100110010000;
			in = 0;
			$monitor("A1 = %b, A2 = %b,in = %b : S = %b,C=%b",A1,A2,in,S,C);
		end



	end
      
endmodule

